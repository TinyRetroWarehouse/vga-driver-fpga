module kord_logo_lut (
	input [9:0] x_i,
	input [8:0] y_i,
	output red_o,
	output green_o,
	output blue_o
);

reg red;
reg green;
reg blue;

assign red_o = red;
assign green_o = green;
assign blue_o = blue;

always @(*) begin
	red = 1'b0;
	green = 1'b0;
	blue = 1'b0;

	if (y_i == 9'd186)
	begin
		if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd187)
	begin
		if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd188)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd189)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd190)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd191)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd192)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd193)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd194)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd195)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd196)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd197)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd198)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd199)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd200)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd201)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd202)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd203)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd204)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd205)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd206)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd207)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd208)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd209)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd210)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd211)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd212)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd213)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd214)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd215)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd348)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd216)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd348)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd217)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd348)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd218)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd348)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd219)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd220)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd221)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd222)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd223)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd224)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd345)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd225)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd226)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd337)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd338)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd339)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd340)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd341)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd344)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd227)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd342)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd343)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd228)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd323)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd229)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd230)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd231)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd232)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd233)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd234)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd235)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd236)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd237)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd238)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd239)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd297)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd240)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd297)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd241)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd297)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd242)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd297)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd243)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd297)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd244)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd297)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd245)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd246)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd247)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd248)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd249)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd250)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd296)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd251)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd252)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd253)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd295)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd254)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd255)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd294)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd256)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd257)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd293)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd258)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd238)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd259)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd239)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd260)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd261)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd240)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd262)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd263)
	begin
		 if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd264)
	begin
		 if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd265)
	begin
		 if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd266)
	begin
		 if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd267)
	begin
		 if (x_i == 10'd182)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd361)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd268)
	begin
		 if (x_i == 10'd181)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd362)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd269)
	begin
		 if (x_i == 10'd180)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd278)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd363)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd364)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd270)
	begin
		 if (x_i == 10'd180)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd224)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd225)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd226)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd227)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd228)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd229)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd230)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd231)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd232)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd233)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd234)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd235)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd236)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd237)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd254)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd255)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd256)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd275)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd276)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd277)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd314)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd315)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd316)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd317)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd318)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd319)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd320)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd321)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd322)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd365)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd366)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd367)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd385)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd401)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd402)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd403)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd404)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd405)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd406)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd407)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd408)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd271)
	begin
		 if (x_i == 10'd179)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd193)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd194)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd257)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd258)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd259)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd260)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd261)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd271)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd272)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd273)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd274)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd368)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd369)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd380)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd381)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd382)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd383)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd384)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd272)
	begin
		 if (x_i == 10'd178)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd191)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd192)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd195)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd379)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd273)
	begin
		 if (x_i == 10'd177)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd189)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd190)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd196)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd197)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
	end
	else if (y_i == 9'd274)
	begin
		 if (x_i == 10'd176)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd186)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd187)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd188)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd198)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
	end
	else if (y_i == 9'd275)
	begin
		 if (x_i == 10'd175)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd176)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd184)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd185)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd199)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd200)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
	end
	else if (y_i == 9'd276)
	begin
		 if (x_i == 10'd175)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd176)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd182)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd183)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd201)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
	end
	else if (y_i == 9'd277)
	begin
		 if (x_i == 10'd174)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd175)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd176)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd181)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd202)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
	end
	else if (y_i == 9'd278)
	begin
		 if (x_i == 10'd173)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd174)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd175)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd176)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd179)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd180)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd203)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
	end
	else if (y_i == 9'd279)
	begin
		 if (x_i == 10'd172)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd173)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd174)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd175)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd176)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd177)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd178)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd204)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd414)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd415)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd416)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd417)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd418)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd419)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd420)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd446)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd447)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd448)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd449)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd450)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd451)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd452)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd463)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd464)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd465)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd466)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd467)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd280)
	begin
		 if (x_i == 10'd172)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd173)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd174)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd175)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd176)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd205)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd241)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd242)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd243)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd244)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd245)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd249)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd250)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd251)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd252)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd253)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd412)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd413)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd414)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd415)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd416)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd417)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd418)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd419)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd420)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd421)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd446)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd447)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd448)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd449)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd450)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd451)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd462)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd463)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd464)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd465)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd466)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd467)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd468)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd281)
	begin
		 if (x_i == 10'd171)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd172)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd173)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd174)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd206)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd207)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd348)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd411)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd412)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd413)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd414)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd420)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd421)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd461)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd462)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd463)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd467)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd468)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd282)
	begin
		 if (x_i == 10'd170)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd171)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd208)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd209)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd348)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd411)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd412)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd461)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd462)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd463)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd283)
	begin
		 if (x_i == 10'd209)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd210)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd211)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd326)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd348)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd411)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd412)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd461)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd462)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd463)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd284)
	begin
		 if (x_i == 10'd211)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd212)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd327)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd411)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd462)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd463)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd464)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd285)
	begin
		 if (x_i == 10'd212)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd213)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd304)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd328)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd411)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd446)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd447)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd448)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd449)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd450)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd451)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd463)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd464)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd465)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd466)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd286)
	begin
		 if (x_i == 10'd213)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd214)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd304)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd305)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd306)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd307)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd308)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd309)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd310)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd329)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd411)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd417)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd418)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd419)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd420)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd421)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd446)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd447)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd448)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd449)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd450)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd451)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd464)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd465)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd466)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd467)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd287)
	begin
		 if (x_i == 10'd214)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd215)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd216)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd279)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd311)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd330)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd409)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd411)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd417)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd418)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd419)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd420)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd421)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd465)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd466)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd467)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd468)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd288)
	begin
		 if (x_i == 10'd216)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd217)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd331)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd346)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd348)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd360)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd386)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd400)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd411)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd420)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd421)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd467)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd468)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd289)
	begin
		 if (x_i == 10'd217)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd218)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd219)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd280)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd348)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd410)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd411)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd412)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd420)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd421)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd467)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd468)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd290)
	begin
		 if (x_i == 10'd219)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd220)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd281)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd332)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd347)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd348)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd359)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd387)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd399)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd411)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd412)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd413)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd420)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd421)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd461)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd462)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd467)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd468)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd291)
	begin
		 if (x_i == 10'd220)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd221)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd282)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd292)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd333)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd348)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd357)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd358)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd388)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd389)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd397)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd398)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd412)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd413)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd414)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd415)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd416)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd417)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd418)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd419)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd420)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd421)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd446)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd447)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd448)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd449)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd450)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd451)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd461)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd462)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd463)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd464)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd465)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd466)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd467)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd468)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd292)
	begin
		 if (x_i == 10'd221)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd222)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd223)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd246)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd247)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd248)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd262)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd263)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd264)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd265)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd266)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd267)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd268)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd269)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd270)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd283)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd284)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd285)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd288)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd289)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd290)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd291)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd301)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd302)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd303)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd312)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd313)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd324)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd325)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd334)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd335)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd336)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd349)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd350)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd351)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd355)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd356)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd370)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd371)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd372)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd373)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd374)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd375)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd376)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd377)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd378)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd390)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd391)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd392)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd395)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd396)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd413)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd414)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd415)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd416)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd417)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd418)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd419)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd420)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd421)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd432)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd433)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd444)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd445)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd446)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd447)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd448)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd449)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd450)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd451)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd452)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd462)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd463)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd464)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd465)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd466)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd467)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
	else if (y_i == 9'd293)
	begin
		if (x_i == 10'd223)
		begin
			red = 1'b0;
			green = 1'b1;
			blue = 1'b0;
		end
		else if (x_i == 10'd286)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd287)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd352)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd353)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd354)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd393)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd394)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd416)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd417)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd418)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd464)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
		else if (x_i == 10'd465)
		begin
			red = 1'b1;
			green = 1'b1;
			blue = 1'b1;
		end
	end
end

endmodule
